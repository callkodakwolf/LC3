package decode_pkg;
	`define BR    4'b0000;
	`define JMP   4'b1100;
	`define ADD   4'b0001;
	`define AND   4'b0101;
	`define NOT   4'b1001;
	`define LD    4'b0010;
	`define LDR    4'b0110;
	`define LDI    4'b1010;
	`define LEA    4'b1110;
	`define ST    4'b0011;
	`define STR    4'b0111:
	`define STI    4'b1011;
endpackage 
