
module memory_access(
						input clk,
						input rst,
						inpit